<?xml version="1.0" encoding="utf-8"?>
<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML 1.0 Transitional//EN" "http://www.w3.org/TR/xhtml1/DTD/xhtml1-transitional.dtd">
<html xmlns="http://www.w3.org/1999/xhtml" xml:lang="sv" lang="sv"><head>
<meta http-equiv="content-type" content="text/html; charset=UTF-8" />



  <title>Hj&auml;lpsida f&ouml;r presentationer</title><style type="text/css"><!-- 
     body {
        font-family: sans-serif;
        margin: 10%;
     }
     .copyright { font-size: smaller } -->
  </style>
  <script type="text/javascript"><!--
    window.onload = load;
    function load()
    {
      var back = document.getElementById("back");
      back.focus();
    }
    // -->  </script>
</head><body>
<h1>Hj&auml;lpsida f&ouml;r presentationer</h1>

<p align="justify">Denna presentation kan anv&auml;ndas p&aring; liknande s&auml;tt som Power Point.
F&ouml;r att bl&auml;ddra till n&auml;sta sida g&aring;r det att trycka p&aring; mellanslagstangenten eller klicka med musens
v&auml;stra knapp s&aring; gott som var som helst p&aring; sidan. Bl&auml;ddra fram&aring;t och
bak&aring;t med h&ouml;ger- respektive v&auml;nsterpiltangenterna eller tangenterna &raquo;Pg&nbsp;Dn&raquo; respektive
&raquo;Pg&nbsp;Up&raquo;. Textens storlek anpassas automatiskt efter webbl&auml;sarens
f&ouml;nsterbredd, men den g&aring;r &auml;ven att justera manuellt med
tangenterna &raquo;S&raquo; och &raquo;B&raquo; f&ouml;r att f&ouml;rminska respektive f&ouml;rstora texten. Alternativt kan
tangenterna &raquo;&lt;&raquo; respektive &raquo;&gt;&raquo; anv&auml;ndas. Tangenten
&raquo;F&raquo; anv&auml;nds f&ouml;r att visa&nbsp;/ d&ouml;lja statusraden l&auml;ngst ner i f&ouml;nstret. Tangenten &raquo;K&raquo;
kopplar p&aring;&nbsp;/ av m&ouml;jligheten att klicka med musen f&ouml;r att bl&auml;ddra till n&auml;sta sida. Tangenten
&raquo;C&raquo; anv&auml;nds f&ouml;r att visa inneh&aring;llsf&ouml;rteckningen och en tryckning p&aring; vilken annan tangent som
helst d&ouml;ljer den. En tryckning p&aring; tangenten &raquo;H&raquo; visar denna hj&auml;lpsida. Tangenten &raquo;F11&raquo;
v&auml;xlar mellan fullsk&auml;rmsvisning och visning i webbl&auml;sarens f&ouml;nster. Observera att vissa webbl&auml;sare kan
ha reserverat n&aring;gra av dessa tangenttryckningar f&ouml;r andra funktioner; detta varierar mellan olika webbl&auml;sare.</p>

<p align="justify"><span lang="en">Firefox</span>anv&auml;ndare kan vid behov installera <a href="http://www.krickelkrackel.de/autohide" lang="en" hreflang="en">autohide</a>
f&ouml;r att verktygsf&auml;lten skall d&ouml;ljas vid &ouml;verg&aring;ng till fullsk&auml;rmsvisning med F11.</p>

<p align="justify">F&ouml;r att se hur <em lang="en">Slidy</em> fungerar, titta p&aring; XHTML-koden genom att v&auml;lja &raquo;Visa
k&auml;lla&raquo; (eller liknande) i webbl&auml;sarens meny eller l&auml;s f&ouml;ljande <a href="http://www.w3.org/Talks/Tools/Slidy/">l&auml;ngre
beskrivning</a>, d&auml;r &auml;ven ytterligare finesser beskrivs. Varje sida &auml;r markerad som
<span lang="en">div</span>-element med attributet <code lang="en">class=&quot;slide&quot;</code>. CSS-positionering och procentuell bredd
kan anv&auml;ndas f&ouml;r att placera bilderna i r&auml;tt skala i f&ouml;rh&aring;llande till
webbl&auml;sarens f&ouml;nsterstorlek. Det som skall visas inkrementiellt
markeras med <code lang="en">class=&quot;incremental&quot;</code>. L&auml;nkar h&auml;nvisar till n&aring;gra skript och stilmallar
som har testats med en m&auml;ngd nutida webbl&auml;sare och bildar ett webbaserat alternativ till propriet&auml;ra
presentationsprogram. St&ouml;d f&ouml;r integrerad editering h&aring;ller p&aring; att utvecklas. Skicka g&auml;rna
kommentarer till <a href="http://www.w3.org/People/Raggett/" lang="en" hreflang="en">Dave
Raggett</a> &lt;<a href="mailto:dsr@w3.org">dsr@w3.org</a>&gt;.
Om du finner <em lang="en">Slidy</em> anv&auml;ndbar kan du &ouml;verv&auml;ga att bli
<a href="http://www.w3.org/Consortium/sup" lang="en" hreflang="en">W3C Supporter</a>.</p>

<p><em>V&auml;lkommen att anv&auml;nda presentationens stilmallar, skript och hj&auml;lpfiler enligt reglerna
f&ouml;r W3C:s <a href="http://www.w3.org/Consortium/Legal/copyright-documents" lang="en" hreflang="en">document use</a>
och <a href="http://www.w3.org/Consortium/Legal/copyright-software" lang="en" hreflang="en">software
licensing</a>!</em></p>

<button id="back" onclick="history.go(-1)">Tillbaka till presentationen</button>

<hr />

<p class="copyright" lang="en"><a rel="Copyright" href="http://www.w3.org/Consortium/Legal/ipr-notice#Copyright">Copyright</a> &copy; 2005
<a href="http://www.w3.org/" shape="rect"><acronym title="World Wide Web Consortium">W3C</acronym></a><sup>&copy;</sup> (<a href="http://www.csail.mit.edu/"><acronym title="Massachusetts Institute of Technology">MIT</acronym></a>,
<a href="http://www.ercim.org/"><acronym title="European Research Consortium for Informatics and Mathematics">ERCIM</acronym></a>,
<a href="http://www.keio.ac.jp/">Keio</a>), All Rights Reserved. W3C
<a href="http://www.w3.org/Consortium/Legal/ipr-notice#Legal_Disclaimer">liability</a>,
<a href="http://www.w3.org/Consortium/Legal/ipr-notice#W3C_Trademarks">trademark</a>,
<a rel="Copyright" href="http://www.w3.org/Consortium/Legal/copyright-documents">document use</a> and <a rel="Copyright" href="http://www.w3.org/Consortium/Legal/copyright-software">software
licensing</a> rules apply.</p>
</body></html>
